netcdf isomip_ice_shelf1 {
dimensions:
	ny = 240 ;
	nx = 40 ;
variables:
	double thick(ny, nx) ;
		thick:units = "m" ;
		thick:standard_name = "ice shelf thickness" ;
	double area(ny, nx) ;
		area:units = "m2" ;
		area:standard_name = "ice shelf area" ;
}
